// A simple AND function
module simple_and(f,x,y);
    input x,y;
    output f;
    assign f= (x&y);
endmodule